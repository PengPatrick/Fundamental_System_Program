module WTM(A, B, Prod, Cout);
	input [3:0] A;
	input [3:0] B;
	output Prod;
	output Cout;



endmodule
