module Mux_32b_8to1(in0, in1, in2, in3, in4, in5, in6, in7, sel, Out);
	
	input [31:0] in0, in1, in2, in3, in4, in5, in6, in7;
	input [2:0] sel;
	output [31:0] Out;
	
	wire [31:0] first, second;
	
	Mux_32b_4to1 mux41(in0, in1, in2, in3, sel[1:0], first);
	Mux_32b_4to1 mux42(in4, in5, in6, in7, sel[1:0], second);
	Mux_32b_2to1 mux21(first, second, sel[2], Out);

endmodule
